
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.config.all;

entity memory_stage is
port(
    rst, clk:IN std_logic;

    stack_in: IN std_logic_vector(1 downto 0);

    writeback_in, ldm_in, port_read_in, mem_to_reg_in: IN std_logic;
    pc_to_stack_in, mem_read_in, mem_write_in, rti_in, ret_in, call_in: IN std_logic;
    int_in: In std_logic_vector(1 downto 0);
    addr_Rsrc1_in, addr_Rsrc2_in, addr_Rdst_in: IN std_logic_vector(2 downto 0);

    alu_result_in, immediate_value_in, rsrc1_data_in: IN std_logic_vector(15 downto 0);
    pc_in: IN std_logic_vector(31 downto 0);

    empty_sp_exception_out, invalid_address_exception_out: OUT std_logic;
    writeback_out, ldm_out, port_read_out, mem_to_reg_out: OUT std_logic;

    addr_Rsrc1_out, addr_Rsrc2_out, addr_Rdst_out: OUT std_logic_vector(2 downto 0);

    memory_data_out: OUT std_logic_vector(31 downto 0);
    alu_result_out, immediate_value_out: OUT std_logic_vector(15 downto 0);
    pc_out: OUT std_logic_vector(31 downto 0)

);
end entity memory_stage;

architecture memory_imp1 of memory_stage is
signal sp: std_logic_vector(31 downto 0);
signal mux_chosen_data_in: std_logic_vector(31 downto 0);
signal mux_chosen_address: std_logic_vector(ADDRESS_SIZE downto 0); --address size
signal can_mem_write, can_mem_read, invalid_address_exception, empty_sp_exception: std_logic;

begin
    -- Update the stack pointer. Falling edge triggered
    update_sp: entity work.update_stack port map(rst, sp, stack_in, int_in, clk, call_in, rti_in, ret_in, sp);
    
    --Exception Triggers [combinational]
    check_sp_exception: entity work.sp_exception_checker port map(sp, stack_in, clk, rti_in, ret_in, empty_sp_exception);
    address_checker_lavel: entity work.address_checker port map(alu_result_in, mem_read_in, mem_write_in, stack_in, invalid_address_exception);
    invalid_address_exception_out <= invalid_address_exception;
    empty_sp_exception_out <= empty_sp_exception;
    --Note: Address to check would be alu result only, we won't do invalid checking on sp!
    --NOTE: The address checker will check for invalidity when its a real address (i.e when memWrite or memRead is activated) 
    
    data_memory_label: entity work.data_memory port map(
        mux_chosen_data_in, mux_chosen_address,
        clk, pc_to_stack_in, can_mem_read, can_mem_write,
        stack_in, rti_in, ret_in,
        memory_data_out
    );

    --ASK: What read if an invalid address? Xs ?
    can_mem_write <= mem_write_in and (not invalid_address_exception) and (not empty_sp_exception); 
    
    can_mem_read <= mem_read_in  and (not invalid_address_exception) and (not empty_sp_exception);
    -- Mux to chose the data to be stored in memory [pc pushing or store a value]
    mux_chosen_data_in <= pc_in when pc_to_stack_in = '1'
                        else (31 downto 16 => '0') & rsrc1_data_in;
    
    -- Mux to chose the address of memory [sp or offset calculated from alu]
    mux_chosen_address <= (ADDRESS_SIZE downto 16 => '0') & alu_result_in when stack_in = "00"
                        else sp(ADDRESS_SIZE downto 0); --NOTE: some left-bits will be truncated from the sp
    
    -- Transfer to the write back buffer
    writeback_out <= writeback_in;
    ldm_out <= ldm_in;
    port_read_out <= port_read_in;
    mem_to_reg_out <= mem_to_reg_in;
    addr_Rsrc1_out <= addr_Rsrc1_in;
    addr_Rsrc2_out <= addr_Rsrc2_in;
    addr_Rdst_out <= addr_Rdst_in;
    alu_result_out <= alu_result_in;
    immediate_value_out <= immediate_value_in;
    pc_out <= pc_in;
end memory_imp1;